*Negative Differential Resistance

.include DiffAmp.txt

VDD   1  0  5
VSS   2  0 -5

x1    3 4 1 2 5 DIFFAMP

Vin   3 0 sin(0 100m 1k 0 0)
R     3 5 100
R1    4 5 1k
R2    4 0 1k

.tran 5u 1

.control
run

set hcopydevtype = postscript
set hcopypscolor = 1
hardcopy NegDiffRes.ps v(3) vs v(3)/100-v(5)/100

.endc
.end
