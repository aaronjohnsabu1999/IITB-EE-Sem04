*Wien Bridge Oscillator

.include DiffAmp.txt

VDD   1  0  5
VSS   2  0 -5

x1    3 4 1 2 5 DIFFAMP

Ra    3 0 1k
Rb    6 5 1k
Ca    3 0 0.142u
Cb    3 6 0.142u
R1    4 5 2.5k
R2    4 0 1k

.tran 0.1u 110m 100m

.control
run

set hcopydevtype = postscript
set hcopypscolor = 1
hardcopy WienBridgeOscillator.ps v(5)

.endc
.end
