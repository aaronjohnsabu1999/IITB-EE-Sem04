*Low Pass Filter

.include DiffAmp.txt

VDD   1  0  5
VSS   2  0 -5

x1    3 4 1 2 5 DIFFAMP

Vp    3 0 0
Vm    6 0 ac 1 dc 0
R1    4 6 150
R2    4 5 480
C1    4 5 100n

.ac dec 10 1 500k

.control
run

set hcopydevtype = postscript
set hcopypscolor = 1
hardcopy LowPassFilter.ps vdb(5) xlog

.endc
.end
