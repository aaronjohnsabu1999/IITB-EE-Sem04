*Band Pass Filter

.include DiffAmp.txt

VDD   1  0  5
VSS   2  0 -5

x1    3 4 1 2 5 DIFFAMP

Vp    3 0 0
Vm    6 0 ac 1 dc 0
R1    7 6 30
R2    5 4 1Meg
C1    4 7 1n
C2    5 7 100n
R3    5 7 100


.ac dec 10 1 500k

.control
run

set hcopydevtype = postscript
set hcopypscolor = 1
hardcopy BandPassFilter.ps vdb(5) xlog

.endc
.end
